// Code your testbench here
// or browse Examples
`include "milestone2_quicktest_tb.sv"